`include "mycpu.svh"

import mycpu_pkg::*;

program rb_test
  (
   input logic 	       clk,
   input logic 	       rst_n,
   output logic [15:0] d_in,
   output logic        rw_in,
   output logic [11:0] rs_in,
   input logic [15:0]  a_out,
   input logic [15:0]  b_out
   );
`protected
    MTI!#j,ZOBi3w'*wx~R>?'sB!!{$iZouBIZVT=?7ZiN"#a[ik]}[F[#*OGQ^W[,Q!!+^=v@tQAY}
    =H=A+YVa^3I[o;lV$r55]XZEjC!WB{Dkihx?zlj?xB#XrBDX,KUtImQ3Cre-Zo1W5]lr[?~jv>E7
    }ZsQ5JE6$~XGG@},v~O7\#*^C}wlqDQu@N]H+l[D*e&$[2KA+3Vf\|H13lCbf2,#VviOstv@Z_Rs
    R<<jHmwY#@}#n+]OXZDEpxlRWjZTrD/Qrw[R?3@c*3C,N^*\1Fis"}2u}dN^=@~KwJ,+Y@TpRJE_
    *mJee[{Yw+UbER#><1?ePppRiU{}s1ArQ&KIKol}I[.4BkT]gA^mIcaT-2XeJn^}3{x3vRhQb[r3
    U]l#7*RRT?To}wp2#zsT!qE<H;un*p\{\[OF#sCH-aY'^!n'A7*{lG\]rr[rAx25;{A>G{2DZ{YB
    VWJ*5\7{<jriHo#]}+-B<Ei<beIu,'RT=V=YTnp"/;Q5WJV<e*}Rj@Vn53]?~X$m!'JHjOrJB*Cn
    ?ev!Q\1<*OVJ>'Z-w#G#[_\JaBYuUOB{#pABaDQ${nwJu~D*'$C<kzZ\Ox~5De3-AjY@*t[,pA|o
    u[~tvR,jxJ'l6}}w_vX>O_7@2l$~!,ru+N,kBG|\2a\@Hj'@7
`endprotected
endprogram
